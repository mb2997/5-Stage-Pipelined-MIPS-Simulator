package mips_pkg;


endpackage : mips_pkg